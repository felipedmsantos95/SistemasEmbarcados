package felipe is
type estado is (inicial, espera, piscaVerdeVec, luzAmarelaVec, luzVermelhaVec, atravessa, PiscaVerdePed, luzVermelhaPed);
end felipe;