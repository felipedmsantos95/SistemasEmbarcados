package felipe is
type estado is (inicial, espera, piscaVerdeVec, luzAmarelaVec, luzVermelhaVec, atravessa, piscaVerdePed, luzVermelhaPed);
end felipe;