package felipe is
type estado is (inicial, parado, contagem);
end felipe